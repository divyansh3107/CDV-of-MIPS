interface inf;
  
  logic memWrite;
  logic [31:0] address;
  logic [31:0] writedata;
  logic [31:0] readdata;
 
endinterface

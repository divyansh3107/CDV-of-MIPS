interface inf();

logic branch;
logic update;
logic prediction;

endinterface
interface inf();
    //logic clk;

  	logic             			  ctrl;
  	logic [4:0]                   in1;
  	logic [4:0]                   in2;

  	logic [4:0]             	  out;     

//   	initial clk <=0;
//     always #10 clk = ~clk;
  
endinterface
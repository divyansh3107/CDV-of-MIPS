interface inf();
   // logic clk;

  	logic [1:0]            		  ctrl;
  	logic [31:0]                   in1;
  	logic [31:0]                   in2;
  logic [31:0]                   in3;
  logic [31:0]                   in4;
  
  	logic [31:0]             	  out;     

//   	initial clk <=0;
//     always #10 clk = ~clk;
  
endinterface
class driver;
    virtual inf vif;
    event drv_done;
    mailbox drv_mbx;

    task run();
        //$display ("T=%0t [Driver] starting ...", $time);

        forever begin
            Packet tr;
            //$display ("T=%0t [Driver] waiting for item ...", $time);
            drv_mbx.get(tr);
          @(*)
            //tr.print("Driver");
            //vif.clk <= tr.clk;
            vif.instcode <= tr.instcode;
            vif.PCSelectE <= tr.PCSelectE;
            vif.PCSelectD <= tr.PCSelectD;
            vif.regWrite <= tr.regWrite;
            vif.regDst <= tr.regDst;
            vif.memWrite <= tr.memWrite;
            vif.aluSrc <= tr.aluSrc;
            vif.memtoReg <= tr.memtoReg;
            vif.branchD <= tr.branchD;
            vif.ALUcontrolD <= tr.ALUcontrolD;
            ->drv_done;
        end
    endtask
endclass